// sistema.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module sistema (
		output wire [1:0] button_external_connection_export, // button_external_connection.export
		output wire [9:0] buzzer_external_connection_export, // buzzer_external_connection.export
		input  wire       clk_clk,                           //                        clk.clk
		input  wire       reset_reset_n,                     //                      reset.reset_n
		output wire [3:0] svsd0_external_connection_export,  //  svsd0_external_connection.export
		output wire [3:0] svsd1_external_connection_export,  //  svsd1_external_connection.export
		output wire [3:0] svsd2_external_connection_export,  //  svsd2_external_connection.export
		output wire [3:0] svsd3_external_connection_export,  //  svsd3_external_connection.export
		output wire [3:0] svsd4_external_connection_export,  //  svsd4_external_connection.export
		output wire [3:0] svsd5_external_connection_export,  //  svsd5_external_connection.export
		output wire [7:0] switch_external_connection_export  // switch_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [15:0] cpu_data_master_address;                              // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                 // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [15:0] cpu_instruction_master_address;                       // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                          // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:UART_avalon_jtag_slave_chipselect -> UART:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_readdata;    // UART:av_readdata -> mm_interconnect_0:UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_waitrequest; // UART:av_waitrequest -> mm_interconnect_0:UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_avalon_jtag_slave_address;     // mm_interconnect_0:UART_avalon_jtag_slave_address -> UART:av_address
	wire         mm_interconnect_0_uart_avalon_jtag_slave_read;        // mm_interconnect_0:UART_avalon_jtag_slave_read -> UART:av_read_n
	wire         mm_interconnect_0_uart_avalon_jtag_slave_write;       // mm_interconnect_0:UART_avalon_jtag_slave_write -> UART:av_write_n
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:UART_avalon_jtag_slave_writedata -> UART:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                  // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                   // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                     // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                 // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         mm_interconnect_0_button_s1_chipselect;               // mm_interconnect_0:BUTTON_s1_chipselect -> BUTTON:chipselect
	wire  [31:0] mm_interconnect_0_button_s1_readdata;                 // BUTTON:readdata -> mm_interconnect_0:BUTTON_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                  // mm_interconnect_0:BUTTON_s1_address -> BUTTON:address
	wire         mm_interconnect_0_button_s1_write;                    // mm_interconnect_0:BUTTON_s1_write -> BUTTON:write_n
	wire  [31:0] mm_interconnect_0_button_s1_writedata;                // mm_interconnect_0:BUTTON_s1_writedata -> BUTTON:writedata
	wire         mm_interconnect_0_buzzer_s1_chipselect;               // mm_interconnect_0:BUZZER_s1_chipselect -> BUZZER:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_s1_readdata;                 // BUZZER:readdata -> mm_interconnect_0:BUZZER_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_s1_address;                  // mm_interconnect_0:BUZZER_s1_address -> BUZZER:address
	wire         mm_interconnect_0_buzzer_s1_write;                    // mm_interconnect_0:BUZZER_s1_write -> BUZZER:write_n
	wire  [31:0] mm_interconnect_0_buzzer_s1_writedata;                // mm_interconnect_0:BUZZER_s1_writedata -> BUZZER:writedata
	wire         mm_interconnect_0_switch_s1_chipselect;               // mm_interconnect_0:SWITCH_s1_chipselect -> SWITCH:chipselect
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                 // SWITCH:readdata -> mm_interconnect_0:SWITCH_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                  // mm_interconnect_0:SWITCH_s1_address -> SWITCH:address
	wire         mm_interconnect_0_switch_s1_write;                    // mm_interconnect_0:SWITCH_s1_write -> SWITCH:write_n
	wire  [31:0] mm_interconnect_0_switch_s1_writedata;                // mm_interconnect_0:SWITCH_s1_writedata -> SWITCH:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_svsd0_s1_chipselect;                // mm_interconnect_0:SVSD0_s1_chipselect -> SVSD0:chipselect
	wire  [31:0] mm_interconnect_0_svsd0_s1_readdata;                  // SVSD0:readdata -> mm_interconnect_0:SVSD0_s1_readdata
	wire   [1:0] mm_interconnect_0_svsd0_s1_address;                   // mm_interconnect_0:SVSD0_s1_address -> SVSD0:address
	wire         mm_interconnect_0_svsd0_s1_write;                     // mm_interconnect_0:SVSD0_s1_write -> SVSD0:write_n
	wire  [31:0] mm_interconnect_0_svsd0_s1_writedata;                 // mm_interconnect_0:SVSD0_s1_writedata -> SVSD0:writedata
	wire         mm_interconnect_0_svsd1_s1_chipselect;                // mm_interconnect_0:SVSD1_s1_chipselect -> SVSD1:chipselect
	wire  [31:0] mm_interconnect_0_svsd1_s1_readdata;                  // SVSD1:readdata -> mm_interconnect_0:SVSD1_s1_readdata
	wire   [1:0] mm_interconnect_0_svsd1_s1_address;                   // mm_interconnect_0:SVSD1_s1_address -> SVSD1:address
	wire         mm_interconnect_0_svsd1_s1_write;                     // mm_interconnect_0:SVSD1_s1_write -> SVSD1:write_n
	wire  [31:0] mm_interconnect_0_svsd1_s1_writedata;                 // mm_interconnect_0:SVSD1_s1_writedata -> SVSD1:writedata
	wire         mm_interconnect_0_svsd2_s1_chipselect;                // mm_interconnect_0:SVSD2_s1_chipselect -> SVSD2:chipselect
	wire  [31:0] mm_interconnect_0_svsd2_s1_readdata;                  // SVSD2:readdata -> mm_interconnect_0:SVSD2_s1_readdata
	wire   [1:0] mm_interconnect_0_svsd2_s1_address;                   // mm_interconnect_0:SVSD2_s1_address -> SVSD2:address
	wire         mm_interconnect_0_svsd2_s1_write;                     // mm_interconnect_0:SVSD2_s1_write -> SVSD2:write_n
	wire  [31:0] mm_interconnect_0_svsd2_s1_writedata;                 // mm_interconnect_0:SVSD2_s1_writedata -> SVSD2:writedata
	wire         mm_interconnect_0_svsd3_s1_chipselect;                // mm_interconnect_0:SVSD3_s1_chipselect -> SVSD3:chipselect
	wire  [31:0] mm_interconnect_0_svsd3_s1_readdata;                  // SVSD3:readdata -> mm_interconnect_0:SVSD3_s1_readdata
	wire   [1:0] mm_interconnect_0_svsd3_s1_address;                   // mm_interconnect_0:SVSD3_s1_address -> SVSD3:address
	wire         mm_interconnect_0_svsd3_s1_write;                     // mm_interconnect_0:SVSD3_s1_write -> SVSD3:write_n
	wire  [31:0] mm_interconnect_0_svsd3_s1_writedata;                 // mm_interconnect_0:SVSD3_s1_writedata -> SVSD3:writedata
	wire         mm_interconnect_0_svsd4_s1_chipselect;                // mm_interconnect_0:SVSD4_s1_chipselect -> SVSD4:chipselect
	wire  [31:0] mm_interconnect_0_svsd4_s1_readdata;                  // SVSD4:readdata -> mm_interconnect_0:SVSD4_s1_readdata
	wire   [1:0] mm_interconnect_0_svsd4_s1_address;                   // mm_interconnect_0:SVSD4_s1_address -> SVSD4:address
	wire         mm_interconnect_0_svsd4_s1_write;                     // mm_interconnect_0:SVSD4_s1_write -> SVSD4:write_n
	wire  [31:0] mm_interconnect_0_svsd4_s1_writedata;                 // mm_interconnect_0:SVSD4_s1_writedata -> SVSD4:writedata
	wire         mm_interconnect_0_svsd5_s1_chipselect;                // mm_interconnect_0:SVSD5_s1_chipselect -> SVSD5:chipselect
	wire  [31:0] mm_interconnect_0_svsd5_s1_readdata;                  // SVSD5:readdata -> mm_interconnect_0:SVSD5_s1_readdata
	wire   [1:0] mm_interconnect_0_svsd5_s1_address;                   // mm_interconnect_0:SVSD5_s1_address -> SVSD5:address
	wire         mm_interconnect_0_svsd5_s1_write;                     // mm_interconnect_0:SVSD5_s1_write -> SVSD5:write_n
	wire  [31:0] mm_interconnect_0_svsd5_s1_writedata;                 // mm_interconnect_0:SVSD5_s1_writedata -> SVSD5:writedata
	wire         irq_mapper_receiver0_irq;                             // TIMER:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // UART:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [BUTTON:reset_n, BUZZER:reset_n, CPU:reset_n, SVSD0:reset_n, SVSD1:reset_n, SVSD2:reset_n, SVSD3:reset_n, SVSD4:reset_n, SVSD5:reset_n, SWITCH:reset_n, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                        // CPU:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> [RAM:reset, mm_interconnect_0:RAM_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;               // rst_controller_001:reset_req -> RAM:reset_req
	wire         rst_controller_002_reset_out_reset;                   // rst_controller_002:reset_out -> [UART:rst_n, mm_interconnect_0:UART_reset_reset_bridge_in_reset_reset]

	sistema_BUTTON button (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_s1_readdata),   //                    .readdata
		.out_port   (button_external_connection_export)       // external_connection.export
	);

	sistema_BUZZER buzzer (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_external_connection_export)       // external_connection.export
	);

	sistema_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	sistema_RAM ram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),       //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),         //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect),    //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),         //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),      //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),     //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable),    //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	sistema_SVSD0 svsd0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_svsd0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_svsd0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_svsd0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_svsd0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_svsd0_s1_readdata),   //                    .readdata
		.out_port   (svsd0_external_connection_export)       // external_connection.export
	);

	sistema_SVSD0 svsd1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_svsd1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_svsd1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_svsd1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_svsd1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_svsd1_s1_readdata),   //                    .readdata
		.out_port   (svsd1_external_connection_export)       // external_connection.export
	);

	sistema_SVSD0 svsd2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_svsd2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_svsd2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_svsd2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_svsd2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_svsd2_s1_readdata),   //                    .readdata
		.out_port   (svsd2_external_connection_export)       // external_connection.export
	);

	sistema_SVSD0 svsd3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_svsd3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_svsd3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_svsd3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_svsd3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_svsd3_s1_readdata),   //                    .readdata
		.out_port   (svsd3_external_connection_export)       // external_connection.export
	);

	sistema_SVSD0 svsd4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_svsd4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_svsd4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_svsd4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_svsd4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_svsd4_s1_readdata),   //                    .readdata
		.out_port   (svsd4_external_connection_export)       // external_connection.export
	);

	sistema_SVSD0 svsd5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_svsd5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_svsd5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_svsd5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_svsd5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_svsd5_s1_readdata),   //                    .readdata
		.out_port   (svsd5_external_connection_export)       // external_connection.export
	);

	sistema_SWITCH switch (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_switch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_switch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_switch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_switch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_switch_s1_readdata),   //                    .readdata
		.out_port   (switch_external_connection_export)       // external_connection.export
	);

	sistema_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	sistema_UART uart (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	sistema_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                            (clk_clk),                                              //                          CLK_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                       //  CPU_reset_reset_bridge_in_reset.reset
		.RAM_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // RAM_reset1_reset_bridge_in_reset.reset
		.UART_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                   // UART_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                (cpu_data_master_address),                              //                  CPU_data_master.address
		.CPU_data_master_waitrequest            (cpu_data_master_waitrequest),                          //                                 .waitrequest
		.CPU_data_master_byteenable             (cpu_data_master_byteenable),                           //                                 .byteenable
		.CPU_data_master_read                   (cpu_data_master_read),                                 //                                 .read
		.CPU_data_master_readdata               (cpu_data_master_readdata),                             //                                 .readdata
		.CPU_data_master_write                  (cpu_data_master_write),                                //                                 .write
		.CPU_data_master_writedata              (cpu_data_master_writedata),                            //                                 .writedata
		.CPU_data_master_debugaccess            (cpu_data_master_debugaccess),                          //                                 .debugaccess
		.CPU_instruction_master_address         (cpu_instruction_master_address),                       //           CPU_instruction_master.address
		.CPU_instruction_master_waitrequest     (cpu_instruction_master_waitrequest),                   //                                 .waitrequest
		.CPU_instruction_master_read            (cpu_instruction_master_read),                          //                                 .read
		.CPU_instruction_master_readdata        (cpu_instruction_master_readdata),                      //                                 .readdata
		.BUTTON_s1_address                      (mm_interconnect_0_button_s1_address),                  //                        BUTTON_s1.address
		.BUTTON_s1_write                        (mm_interconnect_0_button_s1_write),                    //                                 .write
		.BUTTON_s1_readdata                     (mm_interconnect_0_button_s1_readdata),                 //                                 .readdata
		.BUTTON_s1_writedata                    (mm_interconnect_0_button_s1_writedata),                //                                 .writedata
		.BUTTON_s1_chipselect                   (mm_interconnect_0_button_s1_chipselect),               //                                 .chipselect
		.BUZZER_s1_address                      (mm_interconnect_0_buzzer_s1_address),                  //                        BUZZER_s1.address
		.BUZZER_s1_write                        (mm_interconnect_0_buzzer_s1_write),                    //                                 .write
		.BUZZER_s1_readdata                     (mm_interconnect_0_buzzer_s1_readdata),                 //                                 .readdata
		.BUZZER_s1_writedata                    (mm_interconnect_0_buzzer_s1_writedata),                //                                 .writedata
		.BUZZER_s1_chipselect                   (mm_interconnect_0_buzzer_s1_chipselect),               //                                 .chipselect
		.CPU_debug_mem_slave_address            (mm_interconnect_0_cpu_debug_mem_slave_address),        //              CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write              (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                 .write
		.CPU_debug_mem_slave_read               (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                 .read
		.CPU_debug_mem_slave_readdata           (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                 .readdata
		.CPU_debug_mem_slave_writedata          (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                 .writedata
		.CPU_debug_mem_slave_byteenable         (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                 .byteenable
		.CPU_debug_mem_slave_waitrequest        (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                 .waitrequest
		.CPU_debug_mem_slave_debugaccess        (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                 .debugaccess
		.RAM_s1_address                         (mm_interconnect_0_ram_s1_address),                     //                           RAM_s1.address
		.RAM_s1_write                           (mm_interconnect_0_ram_s1_write),                       //                                 .write
		.RAM_s1_readdata                        (mm_interconnect_0_ram_s1_readdata),                    //                                 .readdata
		.RAM_s1_writedata                       (mm_interconnect_0_ram_s1_writedata),                   //                                 .writedata
		.RAM_s1_byteenable                      (mm_interconnect_0_ram_s1_byteenable),                  //                                 .byteenable
		.RAM_s1_chipselect                      (mm_interconnect_0_ram_s1_chipselect),                  //                                 .chipselect
		.RAM_s1_clken                           (mm_interconnect_0_ram_s1_clken),                       //                                 .clken
		.SVSD0_s1_address                       (mm_interconnect_0_svsd0_s1_address),                   //                         SVSD0_s1.address
		.SVSD0_s1_write                         (mm_interconnect_0_svsd0_s1_write),                     //                                 .write
		.SVSD0_s1_readdata                      (mm_interconnect_0_svsd0_s1_readdata),                  //                                 .readdata
		.SVSD0_s1_writedata                     (mm_interconnect_0_svsd0_s1_writedata),                 //                                 .writedata
		.SVSD0_s1_chipselect                    (mm_interconnect_0_svsd0_s1_chipselect),                //                                 .chipselect
		.SVSD1_s1_address                       (mm_interconnect_0_svsd1_s1_address),                   //                         SVSD1_s1.address
		.SVSD1_s1_write                         (mm_interconnect_0_svsd1_s1_write),                     //                                 .write
		.SVSD1_s1_readdata                      (mm_interconnect_0_svsd1_s1_readdata),                  //                                 .readdata
		.SVSD1_s1_writedata                     (mm_interconnect_0_svsd1_s1_writedata),                 //                                 .writedata
		.SVSD1_s1_chipselect                    (mm_interconnect_0_svsd1_s1_chipselect),                //                                 .chipselect
		.SVSD2_s1_address                       (mm_interconnect_0_svsd2_s1_address),                   //                         SVSD2_s1.address
		.SVSD2_s1_write                         (mm_interconnect_0_svsd2_s1_write),                     //                                 .write
		.SVSD2_s1_readdata                      (mm_interconnect_0_svsd2_s1_readdata),                  //                                 .readdata
		.SVSD2_s1_writedata                     (mm_interconnect_0_svsd2_s1_writedata),                 //                                 .writedata
		.SVSD2_s1_chipselect                    (mm_interconnect_0_svsd2_s1_chipselect),                //                                 .chipselect
		.SVSD3_s1_address                       (mm_interconnect_0_svsd3_s1_address),                   //                         SVSD3_s1.address
		.SVSD3_s1_write                         (mm_interconnect_0_svsd3_s1_write),                     //                                 .write
		.SVSD3_s1_readdata                      (mm_interconnect_0_svsd3_s1_readdata),                  //                                 .readdata
		.SVSD3_s1_writedata                     (mm_interconnect_0_svsd3_s1_writedata),                 //                                 .writedata
		.SVSD3_s1_chipselect                    (mm_interconnect_0_svsd3_s1_chipselect),                //                                 .chipselect
		.SVSD4_s1_address                       (mm_interconnect_0_svsd4_s1_address),                   //                         SVSD4_s1.address
		.SVSD4_s1_write                         (mm_interconnect_0_svsd4_s1_write),                     //                                 .write
		.SVSD4_s1_readdata                      (mm_interconnect_0_svsd4_s1_readdata),                  //                                 .readdata
		.SVSD4_s1_writedata                     (mm_interconnect_0_svsd4_s1_writedata),                 //                                 .writedata
		.SVSD4_s1_chipselect                    (mm_interconnect_0_svsd4_s1_chipselect),                //                                 .chipselect
		.SVSD5_s1_address                       (mm_interconnect_0_svsd5_s1_address),                   //                         SVSD5_s1.address
		.SVSD5_s1_write                         (mm_interconnect_0_svsd5_s1_write),                     //                                 .write
		.SVSD5_s1_readdata                      (mm_interconnect_0_svsd5_s1_readdata),                  //                                 .readdata
		.SVSD5_s1_writedata                     (mm_interconnect_0_svsd5_s1_writedata),                 //                                 .writedata
		.SVSD5_s1_chipselect                    (mm_interconnect_0_svsd5_s1_chipselect),                //                                 .chipselect
		.SWITCH_s1_address                      (mm_interconnect_0_switch_s1_address),                  //                        SWITCH_s1.address
		.SWITCH_s1_write                        (mm_interconnect_0_switch_s1_write),                    //                                 .write
		.SWITCH_s1_readdata                     (mm_interconnect_0_switch_s1_readdata),                 //                                 .readdata
		.SWITCH_s1_writedata                    (mm_interconnect_0_switch_s1_writedata),                //                                 .writedata
		.SWITCH_s1_chipselect                   (mm_interconnect_0_switch_s1_chipselect),               //                                 .chipselect
		.TIMER_s1_address                       (mm_interconnect_0_timer_s1_address),                   //                         TIMER_s1.address
		.TIMER_s1_write                         (mm_interconnect_0_timer_s1_write),                     //                                 .write
		.TIMER_s1_readdata                      (mm_interconnect_0_timer_s1_readdata),                  //                                 .readdata
		.TIMER_s1_writedata                     (mm_interconnect_0_timer_s1_writedata),                 //                                 .writedata
		.TIMER_s1_chipselect                    (mm_interconnect_0_timer_s1_chipselect),                //                                 .chipselect
		.UART_avalon_jtag_slave_address         (mm_interconnect_0_uart_avalon_jtag_slave_address),     //           UART_avalon_jtag_slave.address
		.UART_avalon_jtag_slave_write           (mm_interconnect_0_uart_avalon_jtag_slave_write),       //                                 .write
		.UART_avalon_jtag_slave_read            (mm_interconnect_0_uart_avalon_jtag_slave_read),        //                                 .read
		.UART_avalon_jtag_slave_readdata        (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                                 .readdata
		.UART_avalon_jtag_slave_writedata       (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                                 .writedata
		.UART_avalon_jtag_slave_waitrequest     (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.UART_avalon_jtag_slave_chipselect      (mm_interconnect_0_uart_avalon_jtag_slave_chipselect)   //                                 .chipselect
	);

	sistema_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (cpu_debug_reset_request_reset),          // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
